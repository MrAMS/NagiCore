// typedef byte uint8_t;
// typedef shortint uint16_t;
// typedef int uint32_t;
// typedef longint uint64_t;

`define uint8_t byte unsigned
`define uint16_t shortint unsigned
`define uint32_t int unsigned
`define uint64_t longint unsigned
